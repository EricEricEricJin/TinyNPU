`default_nettype none

module eu_wrapper #(
    
) (
    input wire clk, rst_n,

    // to Avalon MM Read: todo

    // to Control Unit RMIO: todo
);
    
endmodule

`default_nettype wire