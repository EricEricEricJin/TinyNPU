`default_nettype none

module rf_ldst_tb;



endmodule

`default_nettype wire 

