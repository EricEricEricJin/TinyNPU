`default_nettype none

function []

`default_nettype wire 