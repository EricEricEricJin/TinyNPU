// `default_nettype none

// class HPS;
//     ref logic clk;
//     ref logic rst_n;
//     ref logic [31:0] h2f_pio32;

//     function new( ref logic clk, ref logic rst_n, ref logic h2f_pio32 );
//         this.clk = clk;
//         this.rst_n = rst_n;
//         this.h2f_pio32 = h2f_pio32;

//         this.h2f_pio32 = 32'h0;
//     endfunction //new()

//     function void load(logic [31:0] sdram_addr, )

//     endfunction

// endclass //HPS


// `default_nettype wire
// automatically generate testbench