// Load and store vector from / to SDRAM

