// fetch from RD, write back to WD 