`default_nettype none

module mat_reg (
    
);
    
endmodule

`default_nettype wire 